(*MSECM(R) GmbH, http://www.msecm.com, info@msecm.com*)
(*Created 2022-2-23, 18:53:21*)
(*Version MSECM(R) Export Module, 6.2020.703*)
(*Wettkampfstrukturliste*)
FORMAT: Wettkampfdefinitionsliste;6;
ERZEUGER: MSECM(R) Export Module;6.2020.703;info@msecm.com;
VERANSTALTUNG: International Swim Meeting Erlangen 2022;Erlangen;50;AUTOMATISCH;
VERANSTALTUNGSORT: Hannah-Stockbauer-Schwimmhalle;Hartmannstraße 121;91058;Erlangen;GER;+49 9131 8234823;;;
AUSSCHREIBUNGIMNETZ: ;
VERANSTALTER: Turnerbund 1888 Erlangen e.V. Schwimmabteilung;
AUSRICHTER: Turnerbund 1888 Erlangen e.V. Schwimmabteilung;;;;;GER;;;;
MELDEADRESSE: ;;;;GER;;;;
MELDESCHLUSS: 21.03.2022;19:00;
BANKVERBINDUNG: Sparkasse Erlangen;DE97763500000000038216;BYLADEM1ERH;
BESONDERES: ;
NACHWEIS: 01.01.2000;17.03.2001;FW;
ABSCHNITT: 1;26.03.2022;08:00;;09:00;N;
ABSCHNITT: 2;26.03.2022;13:15;;14:15;N;
ABSCHNITT: 3;26.03.2022;18:15;;18:30;N;
ABSCHNITT: 4;27.03.2022;07:30;;08:30;N;
ABSCHNITT: 5;27.03.2022;13:30;;14:30;N;
WETTKAMPF: 1;E;1;1;50;B;GL;W;SW;;;
WETTKAMPF: 2;E;1;1;50;B;GL;M;SW;;;
WETTKAMPF: 3;E;1;1;400;F;GL;W;SW;;;
WETTKAMPF: 4;E;1;1;400;F;GL;M;SW;;;
WETTKAMPF: 5;E;1;1;100;S;GL;W;SW;;;
WETTKAMPF: 6;E;1;1;100;S;GL;M;SW;;;
WETTKAMPF: 7;E;1;1;200;B;GL;W;SW;;;
WETTKAMPF: 8;E;1;1;200;B;GL;M;SW;;;
WETTKAMPF: 9;E;2;1;50;F;GL;W;SW;;;
WETTKAMPF: 10;E;2;1;50;F;GL;M;SW;;;
WETTKAMPF: 11;E;2;1;200;L;GL;W;SW;;;
WETTKAMPF: 12;E;2;1;200;L;GL;M;SW;;;
WETTKAMPF: 13;E;2;1;100;R;GL;W;SW;;;
WETTKAMPF: 14;E;2;1;100;R;GL;M;SW;;;
WETTKAMPF: 15;E;3;1;1500;F;GL;W;SW;;;
WETTKAMPF: 16;E;3;1;1500;F;GL;M;SW;;;
WETTKAMPF: 17;E;3;1;800;F;GL;W;SW;;;
WETTKAMPF: 18;E;3;1;800;F;GL;M;SW;;;
WETTKAMPF: 19;E;4;1;50;R;GL;W;SW;;;
WETTKAMPF: 20;E;4;1;50;R;GL;M;SW;;;
WETTKAMPF: 21;E;4;1;200;F;GL;W;SW;;;
WETTKAMPF: 22;E;4;1;200;F;GL;M;SW;;;
WETTKAMPF: 23;E;4;1;100;B;GL;W;SW;;;
WETTKAMPF: 24;E;4;1;100;B;GL;M;SW;;;
WETTKAMPF: 25;E;4;1;200;S;GL;W;SW;;;
WETTKAMPF: 26;E;4;1;200;S;GL;M;SW;;;
WETTKAMPF: 27;E;5;1;50;S;GL;W;SW;;;
WETTKAMPF: 28;E;5;1;50;S;GL;M;SW;;;
WETTKAMPF: 29;E;5;1;200;R;GL;W;SW;;;
WETTKAMPF: 30;E;5;1;200;R;GL;M;SW;;;
WETTKAMPF: 31;E;5;1;100;F;GL;W;SW;;;
WETTKAMPF: 32;E;5;1;100;F;GL;M;SW;;;
WETTKAMPF: 33;E;5;1;400;L;GL;W;SW;;;
WETTKAMPF: 34;E;5;1;400;L;GL;M;SW;;;
WERTUNG: 1;E;10001;JG;2014;2014;W;Jahrgang 2014;
WERTUNG: 1;E;10002;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 1;E;10003;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 1;E;10004;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 1;E;10005;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 1;E;10006;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 1;E;10007;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 1;E;10008;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 1;E;10009;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 1;E;10010;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 1;E;10011;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 2;E;20001;JG;2014;2014;M;Jahrgang 2014;
WERTUNG: 2;E;20002;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 2;E;20003;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 2;E;20004;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 2;E;20005;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 2;E;20006;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 2;E;20007;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 2;E;20008;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 2;E;20009;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 2;E;20010;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 2;E;20011;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 3;E;30001;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 3;E;30002;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 3;E;30003;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 3;E;30004;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 3;E;30005;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 3;E;30006;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 3;E;30007;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 3;E;30008;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 3;E;30009;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 4;E;40001;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 4;E;40002;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 4;E;40003;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 4;E;40004;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 4;E;40005;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 4;E;40006;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 4;E;40007;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 4;E;40008;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 4;E;40009;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 5;E;50001;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 5;E;50002;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 5;E;50003;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 5;E;50004;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 5;E;50005;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 5;E;50006;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 5;E;50007;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 5;E;50008;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 5;E;50009;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 6;E;60001;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 6;E;60002;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 6;E;60003;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 6;E;60004;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 6;E;60005;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 6;E;60006;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 6;E;60007;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 6;E;60008;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 6;E;60009;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 7;E;70001;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 7;E;70002;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 7;E;70003;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 7;E;70004;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 7;E;70005;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 7;E;70006;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 7;E;70007;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 7;E;70008;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 7;E;70009;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 8;E;80001;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 8;E;80002;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 8;E;80003;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 8;E;80004;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 8;E;80005;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 8;E;80006;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 8;E;80007;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 8;E;80008;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 8;E;80009;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 9;E;90001;JG;2014;2014;W;Jahrgang 2014;
WERTUNG: 9;E;90002;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 9;E;90003;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 9;E;90004;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 9;E;90005;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 9;E;90006;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 9;E;90007;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 9;E;90008;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 9;E;90009;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 9;E;90010;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 9;E;90011;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 10;E;100001;JG;2014;2014;M;Jahrgang 2014;
WERTUNG: 10;E;100002;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 10;E;100003;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 10;E;100004;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 10;E;100005;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 10;E;100006;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 10;E;100007;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 10;E;100008;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 10;E;100009;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 10;E;100010;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 10;E;100011;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 11;E;110001;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 11;E;110002;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 11;E;110003;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 11;E;110004;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 11;E;110005;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 11;E;110006;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 11;E;110007;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 11;E;110008;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 11;E;110009;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 12;E;120001;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 12;E;120002;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 12;E;120003;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 12;E;120004;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 12;E;120005;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 12;E;120006;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 12;E;120007;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 12;E;120008;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 12;E;120009;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 13;E;130001;JG;2014;2014;W;Jahrgang 2014;
WERTUNG: 13;E;130002;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 13;E;130003;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 13;E;130004;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 13;E;130005;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 13;E;130006;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 13;E;130007;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 13;E;130008;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 13;E;130009;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 13;E;130010;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 13;E;130011;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 14;E;140001;JG;2014;2014;M;Jahrgang 2014;
WERTUNG: 14;E;140002;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 14;E;140003;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 14;E;140004;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 14;E;140005;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 14;E;140006;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 14;E;140007;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 14;E;140008;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 14;E;140009;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 14;E;140010;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 14;E;140011;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 15;E;150001;JG;0;2011;W;Jahrgang 2011 und älter;
WERTUNG: 16;E;160001;JG;0;2011;M;Jahrgang 2011 und älter;
WERTUNG: 17;E;170001;JG;0;2011;W;Jahrgang 2011 und älter;
WERTUNG: 18;E;180001;JG;0;2011;M;Jahrgang 2011 und älter;
WERTUNG: 19;E;190001;JG;2014;2014;W;Jahrgang 2014;
WERTUNG: 19;E;190002;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 19;E;190003;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 19;E;190004;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 19;E;190005;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 19;E;190006;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 19;E;190007;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 19;E;190008;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 19;E;190009;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 19;E;190010;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 19;E;190011;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 20;E;200001;JG;2014;2014;M;Jahrgang 2014;
WERTUNG: 20;E;200002;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 20;E;200003;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 20;E;200004;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 20;E;200005;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 20;E;200006;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 20;E;200007;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 20;E;200008;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 20;E;200009;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 20;E;200010;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 20;E;200011;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 21;E;210001;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 21;E;210002;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 21;E;210003;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 21;E;210004;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 21;E;210005;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 21;E;210006;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 21;E;210007;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 21;E;210008;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 21;E;210009;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 21;E;210010;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 22;E;220001;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 22;E;220002;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 22;E;220003;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 22;E;220004;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 22;E;220005;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 22;E;220006;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 22;E;220007;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 22;E;220008;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 22;E;220009;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 22;E;220010;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 23;E;230001;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 23;E;230002;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 23;E;230003;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 23;E;230004;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 23;E;230005;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 23;E;230006;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 23;E;230007;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 23;E;230008;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 23;E;230009;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 23;E;230010;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 24;E;240001;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 24;E;240002;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 24;E;240003;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 24;E;240004;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 24;E;240005;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 24;E;240006;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 24;E;240007;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 24;E;240008;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 24;E;240009;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 24;E;240010;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 25;E;250001;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 25;E;250002;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 25;E;250003;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 25;E;250004;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 25;E;250005;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 25;E;250006;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 25;E;250007;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 25;E;250008;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 26;E;260001;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 26;E;260002;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 26;E;260003;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 26;E;260004;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 26;E;260005;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 26;E;260006;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 26;E;260007;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 26;E;260008;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 27;E;270001;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 27;E;270002;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 27;E;270003;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 27;E;270004;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 27;E;270005;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 27;E;270006;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 27;E;270007;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 27;E;270008;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 27;E;270009;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 27;E;270010;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 28;E;280001;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 28;E;280002;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 28;E;280003;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 28;E;280004;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 28;E;280005;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 28;E;280006;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 28;E;280007;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 28;E;280008;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 28;E;280009;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 28;E;280010;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 29;E;290001;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 29;E;290002;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 29;E;290003;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 29;E;290004;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 29;E;290005;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 29;E;290006;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 29;E;290007;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 29;E;290008;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 29;E;290009;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 29;E;290010;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 30;E;300001;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 30;E;300002;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 30;E;300003;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 30;E;300004;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 30;E;300005;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 30;E;300006;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 30;E;300007;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 30;E;300008;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 30;E;300009;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 30;E;300010;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 31;E;310001;JG;2014;2014;W;Jahrgang 2014;
WERTUNG: 31;E;310002;JG;2013;2013;W;Jahrgang 2013;
WERTUNG: 31;E;310003;JG;2012;2012;W;Jahrgang 2012;
WERTUNG: 31;E;310004;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 31;E;310005;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 31;E;310006;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 31;E;310007;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 31;E;310008;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 31;E;310009;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 31;E;310010;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 31;E;310011;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 32;E;320001;JG;2014;2014;M;Jahrgang 2014;
WERTUNG: 32;E;320002;JG;2013;2013;M;Jahrgang 2013;
WERTUNG: 32;E;320003;JG;2012;2012;M;Jahrgang 2012;
WERTUNG: 32;E;320004;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 32;E;320005;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 32;E;320006;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 32;E;320007;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 32;E;320008;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 32;E;320009;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 32;E;320010;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 32;E;320011;JG;0;2004;M;Jahrgang 2004 und älter;
WERTUNG: 33;E;330001;JG;2011;2011;W;Jahrgang 2011;
WERTUNG: 33;E;330002;JG;2010;2010;W;Jahrgang 2010;
WERTUNG: 33;E;330003;JG;2009;2009;W;Jahrgang 2009;
WERTUNG: 33;E;330004;JG;2008;2008;W;Jahrgang 2008;
WERTUNG: 33;E;330005;JG;2007;2007;W;Jahrgang 2007;
WERTUNG: 33;E;330006;JG;2006;2006;W;Jahrgang 2006;
WERTUNG: 33;E;330007;JG;2005;2005;W;Jahrgang 2005;
WERTUNG: 33;E;330008;JG;0;2004;W;Jahrgang 2004 und älter;
WERTUNG: 34;E;340001;JG;2011;2011;M;Jahrgang 2011;
WERTUNG: 34;E;340002;JG;2010;2010;M;Jahrgang 2010;
WERTUNG: 34;E;340003;JG;2009;2009;M;Jahrgang 2009;
WERTUNG: 34;E;340004;JG;2008;2008;M;Jahrgang 2008;
WERTUNG: 34;E;340005;JG;2007;2007;M;Jahrgang 2007;
WERTUNG: 34;E;340006;JG;2006;2006;M;Jahrgang 2006;
WERTUNG: 34;E;340007;JG;2005;2005;M;Jahrgang 2005;
WERTUNG: 34;E;340008;JG;0;2004;M;Jahrgang 2004 und älter;
MELDEGELD: Wkmeldegeld;7,00;1;
MELDEGELD: Wkmeldegeld;7,00;2;
MELDEGELD: Wkmeldegeld;7,00;3;
MELDEGELD: Wkmeldegeld;7,00;4;
MELDEGELD: Wkmeldegeld;7,00;5;
MELDEGELD: Wkmeldegeld;7,00;6;
MELDEGELD: Wkmeldegeld;7,00;7;
MELDEGELD: Wkmeldegeld;7,00;8;
MELDEGELD: Wkmeldegeld;7,00;9;
MELDEGELD: Wkmeldegeld;7,00;10;
MELDEGELD: Wkmeldegeld;7,00;11;
MELDEGELD: Wkmeldegeld;7,00;12;
MELDEGELD: Wkmeldegeld;7,00;13;
MELDEGELD: Wkmeldegeld;7,00;14;
MELDEGELD: Wkmeldegeld;8,00;15;
MELDEGELD: Wkmeldegeld;8,00;16;
MELDEGELD: Wkmeldegeld;8,00;17;
MELDEGELD: Wkmeldegeld;8,00;18;
MELDEGELD: Wkmeldegeld;7,00;19;
MELDEGELD: Wkmeldegeld;7,00;20;
MELDEGELD: Wkmeldegeld;7,00;21;
MELDEGELD: Wkmeldegeld;7,00;22;
MELDEGELD: Wkmeldegeld;7,00;23;
MELDEGELD: Wkmeldegeld;7,00;24;
MELDEGELD: Wkmeldegeld;7,00;25;
MELDEGELD: Wkmeldegeld;7,00;26;
MELDEGELD: Wkmeldegeld;7,00;27;
MELDEGELD: Wkmeldegeld;7,00;28;
MELDEGELD: Wkmeldegeld;7,00;29;
MELDEGELD: Wkmeldegeld;7,00;30;
MELDEGELD: Wkmeldegeld;7,00;31;
MELDEGELD: Wkmeldegeld;7,00;32;
MELDEGELD: Wkmeldegeld;7,00;33;
MELDEGELD: Wkmeldegeld;7,00;34;
DATEIENDE
